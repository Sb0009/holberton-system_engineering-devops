magic
tech minimum
timestamp 1643401545
<< end >>
